module fme(
	clock,
	reset,
	enable,
	in_0,
	in_1,
	in_2,
	in_3,
	in_4,
	in_5,
	in_6,
	in_7,
	in_8,
	in_9,
	in_10,
	in_11,
	in_12,
	in_13,
	in_14,
	in_15,
	in_16,
	in_17,
	in_18,
	in_19,
	in_20,
	in_21,
	in_22,
	in_23,
	in_24,
	in_25,
	in_26,
	in_27,
	in_28,
	in_29,
	in_30,
	in_31,
	out_0,
	out_1,
	out_2,
	out_3,
	out_4,
	out_5,
	out_6,
	out_7,
	out_8,
	out_9,	
	out_10,
	out_11,
	out_12,
	out_13,
	out_14,
	out_15,
	out_16,
	out_17,
	out_18,
	out_19,
	out_20,
	out_21,
	out_22,
	out_23,
	out_24,
	out_25,
	out_26,
	out_27,
	out_28,
	out_29,
	out_30,
	out_31,
	out_32,
	out_33,
	out_34,
	out_35,
	out_36,
	out_37,
	out_38,
	out_39,
	out_40,
	out_41,
	out_42,
	out_43,
	out_44,
	out_45,
	out_46,
	out_47,
	out_48,
	out_49,
	out_50,
	out_51,
	out_52,
	out_53,
	out_54,
	out_55,
	out_56,
	out_57,
	out_58,
	out_59,
	out_60,
	out_61,
	out_62,
	out_63,
	out_64,
	out_65,
	out_66,
	out_67,
	out_68,
	out_69,
	out_70,
	out_71,
	out_72,
	out_73,
	out_74,
	out_75,
	out_76,
	out_77,
	out_78,
	out_79,
	out_80,
	out_81,
	out_82,
	out_83,
	out_84,
	out_85,
	out_86,
	out_87,
	out_88,
	out_89,
	out_90,
	out_91,
	out_92,
	out_93,
	out_94,
	out_95,
	out_96,
	out_97,
	out_98,
	out_99,
	out_100,
	out_101,
	out_102,
	out_103,
	out_104,
	out_105,
	out_106,
	out_107,
	out_108,
	out_109,	
	out_110,
	out_111,
	out_112,
	out_113,
	out_114,
	out_115,
	out_116,
	out_117,
	out_118,
	out_119,
	out_120,
	out_121,
	out_122,
	out_123,
	out_124,
	out_125,
	out_126,
	out_127,
	out_128,
	out_129,
	out_130,
	out_131,
	out_132,
	out_133,
	out_134,
	out_135,
	out_136,
	out_137,
	out_138,
	out_139,
	out_140,
	out_141,
	out_142,
	out_143,
	out_144,
	out_145,
	out_146,
	out_147,
	out_148,
	out_149,
	out_150,
	out_151,
	out_152,
	out_153,
	out_154,
	out_155,
	out_156,
	out_157,
	out_158,
	out_159,
	out_160,
	out_161,
	done
	);


//--------------------------------- Parametros -----------------------------//
 
 parameter DATA_WIDTH = 8;

 //------------------------------- Portas de Entrada -----------------------------------//

input clock, reset, enable;
input [DATA_WIDTH-1:0] in_0, in_1,in_2,in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17,in_18,in_19,in_20,in_21,in_22,in_23,in_24,in_25,in_26, in_27, in_28, in_29, in_30, in_31;

//--------------------------------- Portas de saida -----------------------------//
output [DATA_WIDTH-1:0] out_0,out_1,out_2,out_3,out_4,out_5,out_6,out_7,out_8,out_9,out_10,out_11,out_12,out_13,out_14,out_15,out_16,out_17,out_18,out_19,out_20,out_21,out_22,out_23,out_24,out_25,out_26,out_27,out_28,out_29,out_30,out_31,out_32,out_33,out_34,out_35,out_36,out_37,out_38,out_39,out_40,out_41,out_42,out_43,out_44,out_45,out_46,out_47,out_48,out_49,out_50,out_51,out_52,out_53;

output [DATA_WIDTH-1:0] out_54,out_55,out_56,out_57,out_58,out_59,out_60,out_61,out_62,out_63,out_64,out_65,out_66,out_67,out_68,out_69,out_70,out_71,out_72,out_73,out_74,out_75,out_76,out_77,out_78,out_79,	out_80,out_81,out_82,out_83,out_84,out_85,out_86,out_87,out_88,out_89,	out_90,out_91,out_92,out_93,out_94,out_95,out_96,out_97,out_98,out_99,out_100,out_101,out_102,out_103,out_104,out_105,out_106,out_107,out_108,out_109,	out_110,out_111,out_112,out_113,out_114,out_115,out_116,out_117,out_118,out_119,out_120,out_121,out_122,out_123,out_124,out_125,out_126,out_127,out_128,out_129,out_130,out_131,out_132,out_133,out_134,out_135,out_136,out_137,out_138,out_139,out_140,out_141,out_142,out_143,out_144,out_145,out_146,out_147,out_148,out_149,out_150,out_151,out_152,out_153,out_154,out_155,out_156,out_157,out_158,out_159,out_160,out_161;

output done;

//--------------------------------- Fios Internos -----------------------------//

wire escrita_finalizada, fase1_finalizada, fase2p3_finalizada, fase3_finalizada, pos_interpolacao_finalizada, reseto, enable_buffer_int,direction_buffer_int, modo_leitura, c0, c1, enable_filtros, enable_buffers, direction_buffer_a, direction_buffer_b, direction_buffer_c, enable_buffer_verticais, enable_buffer_diagonais_a, enable_buffer_diagonais_b,enable_buffer_diagonais_c;

//--------------------------------- Bloco de controle e operativo -----------------------------//

fme_controle  #(DATA_WIDTH) fme_con (clock,reset,enable,escrita_finalizada, fase1_finalizada, fase2p3_finalizada,fase3_finalizada, pos_interpolacao_finalizada,reseto,enable_buffer_int,direction_buffer_int,modo_leitura,c0,c1,enable_filtros,enable_buffers,direction_buffer_a,direction_buffer_b,direction_buffer_c,enable_buffer_verticais,enable_buffer_diagonais_a,enable_buffer_diagonais_b,enable_buffer_diagonais_c,done);
fme_operativo #(DATA_WIDTH) fme_op (clock,reset,in_0,in_1,in_2,in_3,in_4,in_5,in_6,in_7,in_8,in_9,in_10,in_11,in_12,in_13,in_14,in_15,in_16,in_17,in_18,in_19,in_20,in_21,in_22,in_23,in_24,in_25,in_26,in_27,in_28,in_29,in_30,in_31,reseto,enable_buffer_int,direction_buffer_int,modo_leitura,c0,c1,enable_filtros,enable_buffers,direction_buffer_a,direction_buffer_b,direction_buffer_c,enable_buffer_verticais,enable_buffer_diagonais_a,enable_buffer_diagonais_b,enable_buffer_diagonais_c,escrita_finalizada, fase1_finalizada, fase2p3_finalizada,fase3_finalizada, pos_interpolacao_finalizada,out_0,out_1,out_2,out_3,out_4,out_5,out_6,out_7,out_8,out_9,out_10,out_11,out_12,out_13,out_14,out_15,out_16,out_17,out_18,out_19,out_20,out_21,out_22,out_23,out_24,out_25,out_26,out_27,out_28,out_29,out_30,out_31,out_32,out_33,out_34,out_35,out_36,out_37,out_38,out_39,out_40,out_41,out_42,out_43,out_44,out_45,out_46,out_47,out_48,out_49,out_50,out_51,out_52,out_53,out_54,out_55,out_56,out_57,out_58,out_59,out_60,out_61,out_62,out_63,out_64,out_65,out_66,out_67,out_68,out_69,out_70,out_71,out_72,out_73,out_74,out_75,out_76,out_77,out_78,out_79,out_80,out_81,out_82,out_83,out_84,out_85,out_86,out_87,out_88,out_89,out_90,out_91,out_92,out_93,out_94,out_95,out_96,out_97,out_98,out_99,out_100,out_101,out_102,out_103,out_104,out_105,out_106,out_107,out_108,out_109,out_110,out_111,out_112,out_113,out_114,out_115,out_116,out_117,out_118,out_119,out_120,out_121,out_122,out_123,out_124,out_125,out_126,out_127,out_128,out_129,out_130,out_131,out_132,out_133,out_134,out_135,out_136,out_137,out_138,out_139,out_140,out_141,out_142,out_143,out_144,out_145,out_146,out_147,out_148,out_149,out_150,out_151,out_152,out_153,out_154,out_155,out_156,out_157,out_158,out_159,out_160,out_161);

endmodule