//`include "buffer_cell.v" 

module buffer_diagonais(
	clock, 
	reset,
	enable,
	in_0,
	in_1,
	in_2,
	in_3,
	in_4,
	in_5,
	in_6,
	in_7,
	in_8,
	in_9,
	in_10,
	in_11,
	in_12,
	in_13,
	in_14,
	in_15,
	in_16,
	in_17,
	in_18,
	in_19,
	in_20,
	in_21,
	in_22,
	in_23,
	in_24,
	in_25,
	in_26,
	out_0,
	out_1,
	out_2,
	out_3,
	out_4,
	out_5,
	out_6,
	out_7,
	out_8,
	out_9,
	out_10,
	out_11,
	out_12,
	out_13,
	out_14,
	out_15,
	out_16,
	out_17,
	out_18,
	out_19,
	out_20,
	out_21,
	out_22,
	out_23,
	out_24,
	out_25,
	out_26
	);

parameter DATA_WIDTH = 8;
input clock, reset, enable;

input signed [DATA_WIDTH+1:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_18,in_19,in_20,in_21,in_22,in_23,in_24,in_25,in_26;
input signed [DATA_WIDTH+2:0] in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17;
output [DATA_WIDTH-1:0] out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15,out_16,out_17,out_18,out_19,out_20,out_21,out_22,out_23,out_24,out_25,out_26;
wire [DATA_WIDTH-1:0] 
out_of_0_0, out_of_0_1, out_of_0_2, out_of_0_3, out_of_0_4, out_of_0_5, out_of_0_6, out_of_0_7, out_of_0_8, 
out_of_1_0, out_of_1_1, out_of_1_2, out_of_1_3, out_of_1_4, out_of_1_5, out_of_1_6, out_of_1_7, out_of_1_8,  
out_of_2_0, out_of_2_1, out_of_2_2, out_of_2_3, out_of_2_4, out_of_2_5, out_of_2_6, out_of_2_7, out_of_2_8, 
out_of_3_0, out_of_3_1, out_of_3_2, out_of_3_3, out_of_3_4, out_of_3_5, out_of_3_6, out_of_3_7, out_of_3_8,  
out_of_4_0, out_of_4_1, out_of_4_2, out_of_4_3, out_of_4_4, out_of_4_5, out_of_4_6, out_of_4_7, out_of_4_8, 
out_of_5_0, out_of_5_1, out_of_5_2, out_of_5_3, out_of_5_4, out_of_5_5, out_of_5_6, out_of_5_7, out_of_5_8, 
out_of_6_0, out_of_6_1, out_of_6_2, out_of_6_3, out_of_6_4, out_of_6_5, out_of_6_6, out_of_6_7, out_of_6_8, 
out_of_7_0, out_of_7_1, out_of_7_2, out_of_7_3, out_of_7_4, out_of_7_5, out_of_7_6, out_of_7_7, out_of_7_8, 
out_of_8_0, out_of_8_1, out_of_8_2, out_of_8_3, out_of_8_4, out_of_8_5, out_of_8_6, out_of_8_7, out_of_8_8, 
out_of_9_0, out_of_9_1, out_of_9_2, out_of_9_3, out_of_9_4, out_of_9_5, out_of_9_6, out_of_9_7, out_of_9_8, 
out_of_10_0, out_of_10_1, out_of_10_2, out_of_10_3, out_of_10_4, out_of_10_5, out_of_10_6, out_of_10_7, out_of_10_8, 
out_of_11_0, out_of_11_1, out_of_11_2, out_of_11_3, out_of_11_4, out_of_11_5, out_of_11_6, out_of_11_7, out_of_11_8, 
out_of_12_0, out_of_12_1, out_of_12_2, out_of_12_3, out_of_12_4, out_of_12_5, out_of_12_6, out_of_12_7, out_of_12_8, 
out_of_13_0, out_of_13_1, out_of_13_2, out_of_13_3, out_of_13_4, out_of_13_5, out_of_13_6, out_of_13_7, out_of_13_8, 
out_of_14_0, out_of_14_1, out_of_14_2, out_of_14_3, out_of_14_4, out_of_14_5, out_of_14_6, out_of_14_7, out_of_14_8, 
out_of_15_0, out_of_15_1, out_of_15_2, out_of_15_3, out_of_15_4, out_of_15_5, out_of_15_6, out_of_15_7, out_of_15_8, 
out_of_16_0, out_of_16_1, out_of_16_2, out_of_16_3, out_of_16_4, out_of_16_5, out_of_16_6, out_of_16_7, out_of_16_8, 
out_of_17_0, out_of_17_1, out_of_17_2, out_of_17_3, out_of_17_4, out_of_17_5, out_of_17_6, out_of_17_7, out_of_17_8, 
out_of_18_0, out_of_18_1, out_of_18_2, out_of_18_3, out_of_18_4, out_of_18_5, out_of_18_6, out_of_18_7, out_of_18_8, 
out_of_19_0, out_of_19_1, out_of_19_2, out_of_19_3, out_of_19_4, out_of_19_5, out_of_19_6, out_of_19_7, out_of_19_8, 
out_of_20_0, out_of_20_1, out_of_20_2, out_of_20_3, out_of_20_4, out_of_20_5, out_of_20_6, out_of_20_7, out_of_20_8, 
out_of_21_0, out_of_21_1, out_of_21_2, out_of_21_3, out_of_21_4, out_of_21_5, out_of_21_6, out_of_21_7, out_of_21_8, 
out_of_22_0, out_of_22_1, out_of_22_2, out_of_22_3, out_of_22_4, out_of_22_5, out_of_22_6, out_of_22_7, out_of_22_8, 
out_of_23_0, out_of_23_1, out_of_23_2, out_of_23_3, out_of_23_4, out_of_23_5, out_of_23_6, out_of_23_7, out_of_23_8, 
out_of_24_0, out_of_24_1, out_of_24_2, out_of_24_3, out_of_24_4, out_of_24_5, out_of_24_6, out_of_24_7, out_of_24_8, 
out_of_25_0, out_of_25_1, out_of_25_2, out_of_25_3, out_of_25_4, out_of_25_5, out_of_25_6, out_of_25_7, out_of_25_8, 
out_of_26_0, out_of_26_1, out_of_26_2, out_of_26_3, out_of_26_4, out_of_26_5, out_of_26_6, out_of_26_7, out_of_26_8;

reg [DATA_WIDTH-1:0] in_0_8bits,in_1_8bits,in_2_8bits,in_3_8bits,in_4_8bits,in_5_8bits,in_6_8bits,in_7_8bits,in_8_8bits,in_9_8bits,
in_10_8bits,in_11_8bits,in_12_8bits,in_13_8bits,in_14_8bits,in_15_8bits,in_16_8bits,in_17_8bits,in_18_8bits,in_19_8bits,
in_20_8bits,in_21_8bits,in_22_8bits,in_23_8bits,in_24_8bits,in_25_8bits,in_26_8bits;


always @ (posedge clock) begin
	if (in_0[9] == 1'b1 ) begin
	in_0_8bits <= 8'b0;
	end else if (in_0[9] == 1'b0 && in_0[8] == 1'b1) begin
  	in_0_8bits <= 8'b11111111;
  	end else begin
	in_0_8bits <= in_0[7:0];
  	end

  	if (in_1[9] == 1'b1 ) begin
	in_1_8bits <= 0;
	end else if (in_1[9] == 1'b0 && in_1[8] == 1'b1) begin
  	in_1_8bits <= 8'b11111111;
  	end else begin
	in_1_8bits <= in_1[7:0];
  	end

  	if (in_2[9] == 1'b1 ) begin
	in_2_8bits <= 0;
	end else if (in_2[9] == 1'b0 && in_2[8] == 1'b1) begin
  	in_2_8bits <= 8'b11111111;
  	end else begin
	in_2_8bits <= in_2[7:0];
  	end

  	if (in_3[9] == 1'b1 ) begin
	in_3_8bits <= 0;
	end else if (in_3[9] == 1'b0 && in_3[8] == 1'b1) begin
  	in_3_8bits <= 8'b11111111;
  	end else begin
	in_3_8bits <= in_3[7:0];
  	end

  	if (in_4[9] == 1'b1 ) begin
	in_4_8bits <= 0;
	end else if (in_4[9] == 1'b0 && in_4[8] == 1'b1) begin
  	in_4_8bits <= 8'b11111111;
  	end else begin
	in_4_8bits <= in_4[7:0];
  	end

  	if (in_5[9] == 1'b1 ) begin
	in_5_8bits <= 0;
	end else if (in_5[9] == 1'b0 && in_5[8] == 1'b1) begin
  	in_5_8bits <= 8'b11111111;
  	end else begin
	in_5_8bits <= in_5[7:0];
  	end

  	if (in_6[9] == 1'b1 ) begin
	in_6_8bits <= 0;
	end else if (in_6[9] == 1'b0 && in_6[8] == 1'b1) begin
  	in_6_8bits <= 8'b11111111;
  	end else begin
	in_6_8bits <= in_6[7:0];
  	end

  	if (in_7[9] == 1'b1 ) begin
	in_7_8bits <= 0;
	end else if (in_7[9] == 1'b0 && in_7[8] == 1'b1) begin
  	in_7_8bits <= 8'b11111111;
  	end else begin
	in_7_8bits <= in_7[7:0];
  	end

  	if (in_8[9] == 1'b1 ) begin
	in_8_8bits <= 0;
	end else if (in_8[9] == 1'b0 && in_8[8] == 1'b1) begin
  	in_8_8bits <= 8'b11111111;
  	end else begin
	in_8_8bits <= in_8[7:0];
  	end

  	if (in_9[10] == 1'b1 ) begin
	in_9_8bits <= 0;
	end else if (in_9[10] == 1'b0 && in_9[8] == 1'b1) begin
  	in_9_8bits <= 8'b11111111;
  	end else begin
	in_9_8bits <= in_9[7:0];
  	end

  	if (in_10[10] == 1'b1 ) begin
	in_10_8bits <= 0;
	end else if (in_10[10] == 1'b0 && in_10[8] == 1'b1) begin
  	in_10_8bits <= 8'b11111111;
  	end else begin
	in_10_8bits <= in_10[7:0];
  	end

  	if (in_11[10] == 1'b1 ) begin
	in_11_8bits <= 0;
	end else if (in_11[10] == 1'b0 && in_11[8] == 1'b1) begin
  	in_11_8bits <= 8'b11111111;
  	end else begin
	in_11_8bits <= in_11[7:0];
  	end

  	if (in_12[10] == 1'b1 ) begin
	in_12_8bits <= 0;
	end else if (in_12[10] == 1'b0 && in_12[8] == 1'b1) begin
  	in_12_8bits <= 8'b11111111;
  	end else begin
	in_12_8bits <= in_12[7:0];
  	end

  	if (in_13[10] == 1'b1 ) begin
	in_13_8bits <= 0;
	end else if (in_13[10] == 1'b0 && in_13[8] == 1'b1) begin
  	in_13_8bits <= 8'b11111111;
  	end else begin
	in_13_8bits <= in_13[7:0];
  	end

  	if (in_14[10] == 1'b1 ) begin
	in_14_8bits <= 0;
	end else if (in_14[10] == 1'b0 && in_14[8] == 1'b1) begin
  	in_14_8bits <= 8'b11111111;
  	end else begin
	in_14_8bits <= in_14[7:0];
  	end

  	if (in_15[10] == 1'b1 ) begin
	in_15_8bits <= 0;
	end else if (in_15[10] == 1'b0 && in_15[8] == 1'b1) begin
  	in_15_8bits <= 8'b11111111;
  	end else begin
	in_15_8bits <= in_15[7:0];
  	end

  	if (in_16[10] == 1'b1 ) begin
	in_16_8bits <= 0;
	end else if (in_16[10] == 1'b0 && in_16[8] == 1'b1) begin
  	in_16_8bits <= 8'b11111111;
  	end else begin
	in_16_8bits <= in_16[7:0];
  	end

  	if (in_17[10] == 1'b1 ) begin
	in_17_8bits <= 0;
	end else if (in_17[10] == 1'b0 && in_17[8] == 1'b1) begin
  	in_17_8bits <= 8'b11111111;
  	end else begin
	in_17_8bits <= in_17[7:0];
  	end

  	if (in_18[9] == 1'b1 ) begin
	in_18_8bits <= 0;
	end else if (in_18[9] == 1'b0 && in_18[8] == 1'b1) begin
  	in_18_8bits <= 8'b11111111;
  	end else begin
	in_18_8bits <= in_18[7:0];
  	end

  	if (in_19[9] == 1'b1 ) begin
	in_19_8bits <= 0;
	end else if (in_19[9] == 1'b0 && in_19[8] == 1'b1) begin
  	in_19_8bits <= 8'b11111111;
  	end else begin
	in_19_8bits <= in_19[7:0];
  	end

  	if (in_20[9] == 1'b1 ) begin
	in_20_8bits <= 0;
	end else if (in_20[9] == 1'b0 && in_20[8] == 1'b1) begin
  	in_20_8bits <= 8'b11111111;
  	end else begin
	in_20_8bits <= in_20[7:0];
  	end

  	if (in_21[9] == 1'b1 ) begin
	in_21_8bits <= 0;
	end else if (in_21[9] == 1'b0 && in_21[8] == 1'b1) begin
  	in_21_8bits <= 8'b11111111;
  	end else begin
	in_21_8bits <= in_21[7:0];
  	end

  	if (in_22[9] == 1'b1 ) begin
	in_22_8bits <= 0;
	end else if (in_22[9] == 1'b0 && in_22[8] == 1'b1) begin
  	in_22_8bits <= 8'b11111111;
  	end else begin
	in_22_8bits <= in_22[7:0];
  	end

  	if (in_23[9] == 1'b1 ) begin
	in_23_8bits <= 0;
	end else if (in_23[9] == 1'b0 && in_23[8] == 1'b1) begin
  	in_23_8bits <= 8'b11111111;
  	end else begin
	in_23_8bits <= in_23[7:0];
  	end

  	if (in_24[9] == 1'b1 ) begin
	in_24_8bits <= 0;
	end else if (in_24[9] == 1'b0 && in_24[8] == 1'b1) begin
  	in_24_8bits <= 8'b11111111;
  	end else begin
	in_24_8bits <= in_24[7:0];
  	end

  	if (in_25[9] == 1'b1 ) begin
	in_25_8bits <= 0;
	end else if (in_25[9] == 1'b0 && in_25[8] == 1'b1) begin
  	in_25_8bits <= 8'b11111111;
  	end else begin
	in_25_8bits <= in_25[7:0];
  	end

  	if (in_26[9] == 1'b1 ) begin
	in_26_8bits <= 0;
	end else if (in_26[9] == 1'b0 && in_26[8] == 1'b1) begin
  	in_26_8bits <= 8'b11111111;
  	end else begin
	in_26_8bits <= in_26[7:0];
  	end
end

buffer_cell #(DATA_WIDTH) cell_0_0(clock, reset, enable, in_0_8bits, out_of_0_0);
buffer_cell #(DATA_WIDTH) cell_1_0(clock, reset, enable, in_1_8bits, out_of_1_0);
buffer_cell #(DATA_WIDTH) cell_2_0(clock, reset, enable, in_2_8bits, out_of_2_0);
buffer_cell #(DATA_WIDTH) cell_3_0(clock, reset, enable, in_3_8bits, out_of_3_0);
buffer_cell #(DATA_WIDTH) cell_4_0(clock, reset, enable, in_4_8bits, out_of_4_0);
buffer_cell #(DATA_WIDTH) cell_5_0(clock, reset, enable, in_5_8bits, out_of_5_0);
buffer_cell #(DATA_WIDTH) cell_6_0(clock, reset, enable, in_6_8bits, out_of_6_0);
buffer_cell #(DATA_WIDTH) cell_7_0(clock, reset, enable, in_7_8bits, out_of_7_0);
buffer_cell #(DATA_WIDTH) cell_8_0(clock, reset, enable, in_8_8bits, out_of_8_0);
buffer_cell #(DATA_WIDTH) cell_9_0(clock, reset, enable, in_9_8bits, out_of_9_0);
buffer_cell #(DATA_WIDTH) cell_10_0(clock, reset, enable, in_10_8bits, out_of_10_0);
buffer_cell #(DATA_WIDTH) cell_11_0(clock, reset, enable, in_11_8bits, out_of_11_0);
buffer_cell #(DATA_WIDTH) cell_12_0(clock, reset, enable, in_12_8bits, out_of_12_0);
buffer_cell #(DATA_WIDTH) cell_13_0(clock, reset, enable, in_13_8bits, out_of_13_0);
buffer_cell #(DATA_WIDTH) cell_14_0(clock, reset, enable, in_14_8bits, out_of_14_0);
buffer_cell #(DATA_WIDTH) cell_15_0(clock, reset, enable, in_15_8bits, out_of_15_0);
buffer_cell #(DATA_WIDTH) cell_16_0(clock, reset, enable, in_16_8bits, out_of_16_0);
buffer_cell #(DATA_WIDTH) cell_17_0(clock, reset, enable, in_17_8bits, out_of_17_0);
buffer_cell #(DATA_WIDTH) cell_18_0(clock, reset, enable, in_18_8bits, out_of_18_0);
buffer_cell #(DATA_WIDTH) cell_19_0(clock, reset, enable, in_19_8bits, out_of_19_0);
buffer_cell #(DATA_WIDTH) cell_20_0(clock, reset, enable, in_20_8bits, out_of_20_0);
buffer_cell #(DATA_WIDTH) cell_21_0(clock, reset, enable, in_21_8bits, out_of_21_0);
buffer_cell #(DATA_WIDTH) cell_22_0(clock, reset, enable, in_22_8bits, out_of_22_0);
buffer_cell #(DATA_WIDTH) cell_23_0(clock, reset, enable, in_23_8bits, out_of_23_0);
buffer_cell #(DATA_WIDTH) cell_24_0(clock, reset, enable, in_24_8bits, out_of_24_0);
buffer_cell #(DATA_WIDTH) cell_25_0(clock, reset, enable, in_25_8bits, out_of_25_0);
buffer_cell #(DATA_WIDTH) cell_26_0(clock, reset, enable, in_26_8bits, out_of_26_0);


buffer_cell #(DATA_WIDTH) cell_0_1(clock, reset, enable,  out_of_0_0,   out_of_0_1);
buffer_cell #(DATA_WIDTH) cell_1_1(clock, reset, enable,  out_of_1_0,   out_of_1_1);
buffer_cell #(DATA_WIDTH) cell_2_1(clock, reset, enable,  out_of_2_0,   out_of_2_1);
buffer_cell #(DATA_WIDTH) cell_3_1(clock, reset, enable,  out_of_3_0,   out_of_3_1);
buffer_cell #(DATA_WIDTH) cell_4_1(clock, reset, enable,  out_of_4_0,   out_of_4_1);
buffer_cell #(DATA_WIDTH) cell_5_1(clock, reset, enable,  out_of_5_0,   out_of_5_1);
buffer_cell #(DATA_WIDTH) cell_6_1(clock, reset, enable,  out_of_6_0,   out_of_6_1);
buffer_cell #(DATA_WIDTH) cell_7_1(clock, reset, enable,  out_of_7_0,   out_of_7_1);
buffer_cell #(DATA_WIDTH) cell_8_1(clock, reset, enable,  out_of_8_0,   out_of_8_1);
buffer_cell #(DATA_WIDTH) cell_9_1(clock, reset, enable,  out_of_9_0,   out_of_9_1);
buffer_cell #(DATA_WIDTH) cell_10_1(clock, reset, enable, out_of_10_0, out_of_10_1);
buffer_cell #(DATA_WIDTH) cell_11_1(clock, reset, enable, out_of_11_0, out_of_11_1);
buffer_cell #(DATA_WIDTH) cell_12_1(clock, reset, enable, out_of_12_0, out_of_12_1);
buffer_cell #(DATA_WIDTH) cell_13_1(clock, reset, enable, out_of_13_0, out_of_13_1);
buffer_cell #(DATA_WIDTH) cell_14_1(clock, reset, enable, out_of_14_0, out_of_14_1);
buffer_cell #(DATA_WIDTH) cell_15_1(clock, reset, enable, out_of_15_0, out_of_15_1);
buffer_cell #(DATA_WIDTH) cell_16_1(clock, reset, enable, out_of_16_0, out_of_16_1);
buffer_cell #(DATA_WIDTH) cell_17_1(clock, reset, enable, out_of_17_0, out_of_17_1);
buffer_cell #(DATA_WIDTH) cell_18_1(clock, reset, enable, out_of_18_0, out_of_18_1);
buffer_cell #(DATA_WIDTH) cell_19_1(clock, reset, enable, out_of_19_0, out_of_19_1);
buffer_cell #(DATA_WIDTH) cell_20_1(clock, reset, enable, out_of_20_0, out_of_20_1);
buffer_cell #(DATA_WIDTH) cell_21_1(clock, reset, enable, out_of_21_0, out_of_21_1);
buffer_cell #(DATA_WIDTH) cell_22_1(clock, reset, enable, out_of_22_0, out_of_22_1);
buffer_cell #(DATA_WIDTH) cell_23_1(clock, reset, enable, out_of_23_0, out_of_23_1);
buffer_cell #(DATA_WIDTH) cell_24_1(clock, reset, enable, out_of_24_0, out_of_24_1);
buffer_cell #(DATA_WIDTH) cell_25_1(clock, reset, enable, out_of_25_0, out_of_25_1);
buffer_cell #(DATA_WIDTH) cell_26_1(clock, reset, enable, out_of_26_0, out_of_26_1);

buffer_cell #(DATA_WIDTH) cell_0_2(clock, reset, enable,   out_of_0_1,  out_of_0_2);
buffer_cell #(DATA_WIDTH) cell_1_2(clock, reset, enable,   out_of_1_1,  out_of_1_2);
buffer_cell #(DATA_WIDTH) cell_2_2(clock, reset, enable,   out_of_2_1,  out_of_2_2);
buffer_cell #(DATA_WIDTH) cell_3_2(clock, reset, enable,   out_of_3_1,  out_of_3_2);
buffer_cell #(DATA_WIDTH) cell_4_2(clock, reset, enable,   out_of_4_1,  out_of_4_2);
buffer_cell #(DATA_WIDTH) cell_5_2(clock, reset, enable,   out_of_5_1,  out_of_5_2);
buffer_cell #(DATA_WIDTH) cell_6_2(clock, reset, enable,   out_of_6_1,  out_of_6_2);
buffer_cell #(DATA_WIDTH) cell_7_2(clock, reset, enable,   out_of_7_1,  out_of_7_2);
buffer_cell #(DATA_WIDTH) cell_8_2(clock, reset, enable,   out_of_8_1,  out_of_8_2);
buffer_cell #(DATA_WIDTH) cell_9_2(clock, reset, enable,   out_of_9_1,  out_of_9_2);
buffer_cell #(DATA_WIDTH) cell_10_2(clock, reset, enable,  out_of_10_1, out_of_10_2);
buffer_cell #(DATA_WIDTH) cell_11_2(clock, reset, enable, out_of_11_1, out_of_11_2);
buffer_cell #(DATA_WIDTH) cell_12_2(clock, reset, enable, out_of_12_1, out_of_12_2);
buffer_cell #(DATA_WIDTH) cell_13_2(clock, reset, enable, out_of_13_1, out_of_13_2);
buffer_cell #(DATA_WIDTH) cell_14_2(clock, reset, enable, out_of_14_1, out_of_14_2);
buffer_cell #(DATA_WIDTH) cell_15_2(clock, reset, enable, out_of_15_1, out_of_15_2);
buffer_cell #(DATA_WIDTH) cell_16_2(clock, reset, enable, out_of_16_1, out_of_16_2);
buffer_cell #(DATA_WIDTH) cell_17_2(clock, reset, enable, out_of_17_1, out_of_17_2);
buffer_cell #(DATA_WIDTH) cell_18_2(clock, reset, enable, out_of_18_1, out_of_18_2);
buffer_cell #(DATA_WIDTH) cell_19_2(clock, reset, enable, out_of_19_1, out_of_19_2);
buffer_cell #(DATA_WIDTH) cell_20_2(clock, reset, enable, out_of_20_1, out_of_20_2);
buffer_cell #(DATA_WIDTH) cell_21_2(clock, reset, enable, out_of_21_1, out_of_21_2);
buffer_cell #(DATA_WIDTH) cell_22_2(clock, reset, enable, out_of_22_1, out_of_22_2);
buffer_cell #(DATA_WIDTH) cell_23_2(clock, reset, enable, out_of_23_1, out_of_23_2);
buffer_cell #(DATA_WIDTH) cell_24_2(clock, reset, enable, out_of_24_1, out_of_24_2);
buffer_cell #(DATA_WIDTH) cell_25_2(clock, reset, enable, out_of_25_1, out_of_25_2);
buffer_cell #(DATA_WIDTH) cell_26_2(clock, reset, enable, out_of_26_1, out_of_26_2);

buffer_cell #(DATA_WIDTH) cell_0_3(clock, reset, enable,   out_of_0_2,  out_of_0_3);
buffer_cell #(DATA_WIDTH) cell_1_3(clock, reset, enable,   out_of_1_2,  out_of_1_3);
buffer_cell #(DATA_WIDTH) cell_2_3(clock, reset, enable,   out_of_2_2,  out_of_2_3);
buffer_cell #(DATA_WIDTH) cell_3_3(clock, reset, enable,   out_of_3_2,  out_of_3_3);
buffer_cell #(DATA_WIDTH) cell_4_3(clock, reset, enable,   out_of_4_2,  out_of_4_3);
buffer_cell #(DATA_WIDTH) cell_5_3(clock, reset, enable,   out_of_5_2,  out_of_5_3);
buffer_cell #(DATA_WIDTH) cell_6_3(clock, reset, enable,   out_of_6_2,  out_of_6_3);
buffer_cell #(DATA_WIDTH) cell_7_3(clock, reset, enable,   out_of_7_2,  out_of_7_3);
buffer_cell #(DATA_WIDTH) cell_8_3(clock, reset, enable,   out_of_8_2,  out_of_8_3);
buffer_cell #(DATA_WIDTH) cell_9_3(clock, reset, enable,   out_of_9_2,  out_of_9_3);
buffer_cell #(DATA_WIDTH) cell_10_3(clock, reset, enable,  out_of_10_2, out_of_10_3);
buffer_cell #(DATA_WIDTH) cell_11_3(clock, reset, enable, out_of_11_2, out_of_11_3);
buffer_cell #(DATA_WIDTH) cell_12_3(clock, reset, enable, out_of_12_2, out_of_12_3);
buffer_cell #(DATA_WIDTH) cell_13_3(clock, reset, enable, out_of_13_2, out_of_13_3);
buffer_cell #(DATA_WIDTH) cell_14_3(clock, reset, enable, out_of_14_2, out_of_14_3);
buffer_cell #(DATA_WIDTH) cell_15_3(clock, reset, enable, out_of_15_2, out_of_15_3);
buffer_cell #(DATA_WIDTH) cell_16_3(clock, reset, enable, out_of_16_2, out_of_16_3);
buffer_cell #(DATA_WIDTH) cell_17_3(clock, reset, enable, out_of_17_2, out_of_17_3);
buffer_cell #(DATA_WIDTH) cell_18_3(clock, reset, enable, out_of_18_2, out_of_18_3);
buffer_cell #(DATA_WIDTH) cell_19_3(clock, reset, enable, out_of_19_2, out_of_19_3);
buffer_cell #(DATA_WIDTH) cell_20_3(clock, reset, enable, out_of_20_2, out_of_20_3);
buffer_cell #(DATA_WIDTH) cell_21_3(clock, reset, enable, out_of_21_2, out_of_21_3);
buffer_cell #(DATA_WIDTH) cell_22_3(clock, reset, enable, out_of_22_2, out_of_22_3);
buffer_cell #(DATA_WIDTH) cell_23_3(clock, reset, enable, out_of_23_2, out_of_23_3);
buffer_cell #(DATA_WIDTH) cell_24_3(clock, reset, enable, out_of_24_2, out_of_24_3);
buffer_cell #(DATA_WIDTH) cell_25_3(clock, reset, enable, out_of_25_2, out_of_25_3);
buffer_cell #(DATA_WIDTH) cell_26_3(clock, reset, enable, out_of_26_2, out_of_26_3);

buffer_cell #(DATA_WIDTH) cell_0_4(clock, reset, enable,   out_of_0_3,  out_of_0_4);
buffer_cell #(DATA_WIDTH) cell_1_4(clock, reset, enable,   out_of_1_3,  out_of_1_4);
buffer_cell #(DATA_WIDTH) cell_2_4(clock, reset, enable,   out_of_2_3,  out_of_2_4);
buffer_cell #(DATA_WIDTH) cell_3_4(clock, reset, enable,   out_of_3_3,  out_of_3_4);
buffer_cell #(DATA_WIDTH) cell_4_4(clock, reset, enable,   out_of_4_3,  out_of_4_4);
buffer_cell #(DATA_WIDTH) cell_5_4(clock, reset, enable,   out_of_5_3,  out_of_5_4);
buffer_cell #(DATA_WIDTH) cell_6_4(clock, reset, enable,   out_of_6_3,  out_of_6_4);
buffer_cell #(DATA_WIDTH) cell_7_4(clock, reset, enable,   out_of_7_3,  out_of_7_4);
buffer_cell #(DATA_WIDTH) cell_8_4(clock, reset, enable,   out_of_8_3,  out_of_8_4);
buffer_cell #(DATA_WIDTH) cell_9_4(clock, reset, enable,   out_of_9_3,  out_of_9_4);
buffer_cell #(DATA_WIDTH) cell_10_4(clock, reset, enable,  out_of_10_3, out_of_10_4);
buffer_cell #(DATA_WIDTH) cell_11_4(clock, reset, enable, out_of_11_3, out_of_11_4);
buffer_cell #(DATA_WIDTH) cell_12_4(clock, reset, enable, out_of_12_3, out_of_12_4);
buffer_cell #(DATA_WIDTH) cell_13_4(clock, reset, enable, out_of_13_3, out_of_13_4);
buffer_cell #(DATA_WIDTH) cell_14_4(clock, reset, enable, out_of_14_3, out_of_14_4);
buffer_cell #(DATA_WIDTH) cell_15_4(clock, reset, enable, out_of_15_3, out_of_15_4);
buffer_cell #(DATA_WIDTH) cell_16_4(clock, reset, enable, out_of_16_3, out_of_16_4);
buffer_cell #(DATA_WIDTH) cell_17_4(clock, reset, enable, out_of_17_3, out_of_17_4);
buffer_cell #(DATA_WIDTH) cell_18_4(clock, reset, enable, out_of_18_3, out_of_18_4);
buffer_cell #(DATA_WIDTH) cell_19_4(clock, reset, enable, out_of_19_3, out_of_19_4);
buffer_cell #(DATA_WIDTH) cell_20_4(clock, reset, enable, out_of_20_3, out_of_20_4);
buffer_cell #(DATA_WIDTH) cell_21_4(clock, reset, enable, out_of_21_3, out_of_21_4);
buffer_cell #(DATA_WIDTH) cell_22_4(clock, reset, enable, out_of_22_3, out_of_22_4);
buffer_cell #(DATA_WIDTH) cell_23_4(clock, reset, enable, out_of_23_3, out_of_23_4);
buffer_cell #(DATA_WIDTH) cell_24_4(clock, reset, enable, out_of_24_3, out_of_24_4);
buffer_cell #(DATA_WIDTH) cell_25_4(clock, reset, enable, out_of_25_3, out_of_25_4);
buffer_cell #(DATA_WIDTH) cell_26_4(clock, reset, enable, out_of_26_3, out_of_26_4);

buffer_cell #(DATA_WIDTH) cell_0_5(clock, reset, enable,   out_of_0_4,  out_of_0_5);
buffer_cell #(DATA_WIDTH) cell_1_5(clock, reset, enable,   out_of_1_4,  out_of_1_5);
buffer_cell #(DATA_WIDTH) cell_2_5(clock, reset, enable,   out_of_2_4,  out_of_2_5);
buffer_cell #(DATA_WIDTH) cell_3_5(clock, reset, enable,   out_of_3_4,  out_of_3_5);
buffer_cell #(DATA_WIDTH) cell_4_5(clock, reset, enable,   out_of_4_4,  out_of_4_5);
buffer_cell #(DATA_WIDTH) cell_5_5(clock, reset, enable,   out_of_5_4,  out_of_5_5);
buffer_cell #(DATA_WIDTH) cell_6_5(clock, reset, enable,   out_of_6_4,  out_of_6_5);
buffer_cell #(DATA_WIDTH) cell_7_5(clock, reset, enable,   out_of_7_4,  out_of_7_5);
buffer_cell #(DATA_WIDTH) cell_8_5(clock, reset, enable,   out_of_8_4,  out_of_8_5);
buffer_cell #(DATA_WIDTH) cell_9_5(clock, reset, enable,   out_of_9_4,  out_of_9_5);
buffer_cell #(DATA_WIDTH) cell_10_5(clock, reset, enable,  out_of_10_4, out_of_10_5);
buffer_cell #(DATA_WIDTH) cell_11_5(clock, reset, enable, out_of_11_4, out_of_11_5);
buffer_cell #(DATA_WIDTH) cell_12_5(clock, reset, enable, out_of_12_4, out_of_12_5);
buffer_cell #(DATA_WIDTH) cell_13_5(clock, reset, enable, out_of_13_4, out_of_13_5);
buffer_cell #(DATA_WIDTH) cell_14_5(clock, reset, enable, out_of_14_4, out_of_14_5);
buffer_cell #(DATA_WIDTH) cell_15_5(clock, reset, enable, out_of_15_4, out_of_15_5);
buffer_cell #(DATA_WIDTH) cell_16_5(clock, reset, enable, out_of_16_4, out_of_16_5);
buffer_cell #(DATA_WIDTH) cell_17_5(clock, reset, enable, out_of_17_4, out_of_17_5);
buffer_cell #(DATA_WIDTH) cell_18_5(clock, reset, enable, out_of_18_4, out_of_18_5);
buffer_cell #(DATA_WIDTH) cell_19_5(clock, reset, enable, out_of_19_4, out_of_19_5);
buffer_cell #(DATA_WIDTH) cell_20_5(clock, reset, enable, out_of_20_4, out_of_20_5);
buffer_cell #(DATA_WIDTH) cell_21_5(clock, reset, enable, out_of_21_4, out_of_21_5);
buffer_cell #(DATA_WIDTH) cell_22_5(clock, reset, enable, out_of_22_4, out_of_22_5);
buffer_cell #(DATA_WIDTH) cell_23_5(clock, reset, enable, out_of_23_4, out_of_23_5);
buffer_cell #(DATA_WIDTH) cell_24_5(clock, reset, enable, out_of_24_4, out_of_24_5);
buffer_cell #(DATA_WIDTH) cell_25_5(clock, reset, enable, out_of_25_4, out_of_25_5);
buffer_cell #(DATA_WIDTH) cell_26_5(clock, reset, enable, out_of_26_4, out_of_26_5);

buffer_cell #(DATA_WIDTH) cell_0_6(clock, reset, enable,   out_of_0_5,  out_of_0_6);
buffer_cell #(DATA_WIDTH) cell_1_6(clock, reset, enable,   out_of_1_5,  out_of_1_6);
buffer_cell #(DATA_WIDTH) cell_2_6(clock, reset, enable,   out_of_2_5,  out_of_2_6);
buffer_cell #(DATA_WIDTH) cell_3_6(clock, reset, enable,   out_of_3_5,  out_of_3_6);
buffer_cell #(DATA_WIDTH) cell_4_6(clock, reset, enable,   out_of_4_5,  out_of_4_6);
buffer_cell #(DATA_WIDTH) cell_5_6(clock, reset, enable,   out_of_5_5,  out_of_5_6);
buffer_cell #(DATA_WIDTH) cell_6_6(clock, reset, enable,   out_of_6_5,  out_of_6_6);
buffer_cell #(DATA_WIDTH) cell_7_6(clock, reset, enable,   out_of_7_5,  out_of_7_6);
buffer_cell #(DATA_WIDTH) cell_8_6(clock, reset, enable,   out_of_8_5,  out_of_8_6);
buffer_cell #(DATA_WIDTH) cell_9_6(clock, reset, enable,   out_of_9_5,  out_of_9_6);
buffer_cell #(DATA_WIDTH) cell_10_6(clock, reset, enable,  out_of_10_5, out_of_10_6);
buffer_cell #(DATA_WIDTH) cell_11_6(clock, reset, enable, out_of_11_5, out_of_11_6);
buffer_cell #(DATA_WIDTH) cell_12_6(clock, reset, enable, out_of_12_5, out_of_12_6);
buffer_cell #(DATA_WIDTH) cell_13_6(clock, reset, enable, out_of_13_5, out_of_13_6);
buffer_cell #(DATA_WIDTH) cell_14_6(clock, reset, enable, out_of_14_5, out_of_14_6);
buffer_cell #(DATA_WIDTH) cell_15_6(clock, reset, enable, out_of_15_5, out_of_15_6);
buffer_cell #(DATA_WIDTH) cell_16_6(clock, reset, enable, out_of_16_5, out_of_16_6);
buffer_cell #(DATA_WIDTH) cell_17_6(clock, reset, enable, out_of_17_5, out_of_17_6);
buffer_cell #(DATA_WIDTH) cell_18_6(clock, reset, enable, out_of_18_5, out_of_18_6);
buffer_cell #(DATA_WIDTH) cell_19_6(clock, reset, enable, out_of_19_5, out_of_19_6);
buffer_cell #(DATA_WIDTH) cell_20_6(clock, reset, enable, out_of_20_5, out_of_20_6);
buffer_cell #(DATA_WIDTH) cell_21_6(clock, reset, enable, out_of_21_5, out_of_21_6);
buffer_cell #(DATA_WIDTH) cell_22_6(clock, reset, enable, out_of_22_5, out_of_22_6);
buffer_cell #(DATA_WIDTH) cell_23_6(clock, reset, enable, out_of_23_5, out_of_23_6);
buffer_cell #(DATA_WIDTH) cell_24_6(clock, reset, enable, out_of_24_5, out_of_24_6);
buffer_cell #(DATA_WIDTH) cell_25_6(clock, reset, enable, out_of_25_5, out_of_25_6);
buffer_cell #(DATA_WIDTH) cell_26_6(clock, reset, enable, out_of_26_5, out_of_26_6);

buffer_cell #(DATA_WIDTH) cell_0_7(clock, reset, enable,   out_of_0_6,  out_of_0_7);
buffer_cell #(DATA_WIDTH) cell_1_7(clock, reset, enable,   out_of_1_6,  out_of_1_7);
buffer_cell #(DATA_WIDTH) cell_2_7(clock, reset, enable,   out_of_2_6,  out_of_2_7);
buffer_cell #(DATA_WIDTH) cell_3_7(clock, reset, enable,   out_of_3_6,  out_of_3_7);
buffer_cell #(DATA_WIDTH) cell_4_7(clock, reset, enable,   out_of_4_6,  out_of_4_7);
buffer_cell #(DATA_WIDTH) cell_5_7(clock, reset, enable,   out_of_5_6,  out_of_5_7);
buffer_cell #(DATA_WIDTH) cell_6_7(clock, reset, enable,   out_of_6_6,  out_of_6_7);
buffer_cell #(DATA_WIDTH) cell_7_7(clock, reset, enable,   out_of_7_6,  out_of_7_7);
buffer_cell #(DATA_WIDTH) cell_8_7(clock, reset, enable,   out_of_8_6,  out_of_8_7);
buffer_cell #(DATA_WIDTH) cell_9_7(clock, reset, enable,   out_of_9_6,  out_of_9_7);
buffer_cell #(DATA_WIDTH) cell_10_7(clock, reset, enable,  out_of_10_6, out_of_10_7);
buffer_cell #(DATA_WIDTH) cell_11_7(clock, reset, enable, out_of_11_6, out_of_11_7);
buffer_cell #(DATA_WIDTH) cell_12_7(clock, reset, enable, out_of_12_6, out_of_12_7);
buffer_cell #(DATA_WIDTH) cell_13_7(clock, reset, enable, out_of_13_6, out_of_13_7);
buffer_cell #(DATA_WIDTH) cell_14_7(clock, reset, enable, out_of_14_6, out_of_14_7);
buffer_cell #(DATA_WIDTH) cell_15_7(clock, reset, enable, out_of_15_6, out_of_15_7);
buffer_cell #(DATA_WIDTH) cell_16_7(clock, reset, enable, out_of_16_6, out_of_16_7);
buffer_cell #(DATA_WIDTH) cell_17_7(clock, reset, enable, out_of_17_6, out_of_17_7);
buffer_cell #(DATA_WIDTH) cell_18_7(clock, reset, enable, out_of_18_6, out_of_18_7);
buffer_cell #(DATA_WIDTH) cell_19_7(clock, reset, enable, out_of_19_6, out_of_19_7);
buffer_cell #(DATA_WIDTH) cell_20_7(clock, reset, enable, out_of_20_6, out_of_20_7);
buffer_cell #(DATA_WIDTH) cell_21_7(clock, reset, enable, out_of_21_6, out_of_21_7);
buffer_cell #(DATA_WIDTH) cell_22_7(clock, reset, enable, out_of_22_6, out_of_22_7);
buffer_cell #(DATA_WIDTH) cell_23_7(clock, reset, enable, out_of_23_6, out_of_23_7);
buffer_cell #(DATA_WIDTH) cell_24_7(clock, reset, enable, out_of_24_6, out_of_24_7);
buffer_cell #(DATA_WIDTH) cell_25_7(clock, reset, enable, out_of_25_6, out_of_25_7);
buffer_cell #(DATA_WIDTH) cell_26_7(clock, reset, enable, out_of_26_6, out_of_26_7);

buffer_cell #(DATA_WIDTH) cell_0_8(clock, reset, enable,   out_of_0_7,  out_of_0_8);
buffer_cell #(DATA_WIDTH) cell_1_8(clock, reset, enable,   out_of_1_7,  out_of_1_8);
buffer_cell #(DATA_WIDTH) cell_2_8(clock, reset, enable,   out_of_2_7,  out_of_2_8);
buffer_cell #(DATA_WIDTH) cell_3_8(clock, reset, enable,   out_of_3_7,  out_of_3_8);
buffer_cell #(DATA_WIDTH) cell_4_8(clock, reset, enable,   out_of_4_7,  out_of_4_8);
buffer_cell #(DATA_WIDTH) cell_5_8(clock, reset, enable,   out_of_5_7,  out_of_5_8);
buffer_cell #(DATA_WIDTH) cell_6_8(clock, reset, enable,   out_of_6_7,  out_of_6_8);
buffer_cell #(DATA_WIDTH) cell_7_8(clock, reset, enable,   out_of_7_7,  out_of_7_8);
buffer_cell #(DATA_WIDTH) cell_8_8(clock, reset, enable,   out_of_8_7,  out_of_8_8);
buffer_cell #(DATA_WIDTH) cell_9_8(clock, reset, enable,   out_of_9_7,  out_of_9_8);
buffer_cell #(DATA_WIDTH) cell_10_8(clock, reset, enable,  out_of_10_7, out_of_10_8);
buffer_cell #(DATA_WIDTH) cell_11_8(clock, reset, enable, out_of_11_7, out_of_11_8);
buffer_cell #(DATA_WIDTH) cell_12_8(clock, reset, enable, out_of_12_7, out_of_12_8);
buffer_cell #(DATA_WIDTH) cell_13_8(clock, reset, enable, out_of_13_7, out_of_13_8);
buffer_cell #(DATA_WIDTH) cell_14_8(clock, reset, enable, out_of_14_7, out_of_14_8);
buffer_cell #(DATA_WIDTH) cell_15_8(clock, reset, enable, out_of_15_7, out_of_15_8);
buffer_cell #(DATA_WIDTH) cell_16_8(clock, reset, enable, out_of_16_7, out_of_16_8);
buffer_cell #(DATA_WIDTH) cell_17_8(clock, reset, enable, out_of_17_7, out_of_17_8);
buffer_cell #(DATA_WIDTH) cell_18_8(clock, reset, enable, out_of_18_7, out_of_18_8);
buffer_cell #(DATA_WIDTH) cell_19_8(clock, reset, enable, out_of_19_7, out_of_19_8);
buffer_cell #(DATA_WIDTH) cell_20_8(clock, reset, enable, out_of_20_7, out_of_20_8);
buffer_cell #(DATA_WIDTH) cell_21_8(clock, reset, enable, out_of_21_7, out_of_21_8);
buffer_cell #(DATA_WIDTH) cell_22_8(clock, reset, enable, out_of_22_7, out_of_22_8);
buffer_cell #(DATA_WIDTH) cell_23_8(clock, reset, enable, out_of_23_7, out_of_23_8);
buffer_cell #(DATA_WIDTH) cell_24_8(clock, reset, enable, out_of_24_7, out_of_24_8);
buffer_cell #(DATA_WIDTH) cell_25_8(clock, reset, enable, out_of_25_7, out_of_25_8);
buffer_cell #(DATA_WIDTH) cell_26_8(clock, reset, enable, out_of_26_7, out_of_26_8);

assign out_0 = out_of_0_8;
assign out_1 = out_of_1_8;
assign out_2 = out_of_2_8;
assign out_3 = out_of_3_8;
assign out_4 = out_of_4_8;
assign out_5 = out_of_5_8;
assign out_6 = out_of_6_8;
assign out_7 = out_of_7_8;
assign out_8 = out_of_8_8;
assign out_9  = out_of_9_8;
assign out_10 = out_of_10_8;
assign out_11 = out_of_11_8;
assign out_12 = out_of_12_8;
assign out_13 = out_of_13_8;
assign out_14 = out_of_14_8;
assign out_15 = out_of_15_8;
assign out_16 = out_of_16_8;
assign out_17 = out_of_17_8;
assign out_18 = out_of_18_8;
assign out_19 = out_of_19_8;
assign out_20 = out_of_20_8;
assign out_21 = out_of_21_8;
assign out_22 = out_of_22_8;
assign out_23 = out_of_23_8;
assign out_24 = out_of_24_8;
assign out_25 = out_of_25_8;
assign out_26 = out_of_26_8;



endmodule
